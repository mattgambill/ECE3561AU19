LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY regLine IS
	PORT (
		ABUS, BBUS                                  : INOUT std_logic_vector(15 DOWNTO 0);
		Aload, Bload, Adrive, Bdrive, Arsel, Brsel  : IN std_logic
	);
END regLine;

ARCHITECTURE one OF regLine IS

	-- define subcomponents
	COMPONENT busdr IS
		PORT (
		     dr       : IN std_logic;
		     datain   : IN std_logic_vector(15 DOWNTO 0);
   		     dataout  : OUT std_logic_vector(15 DOWNTO 0)
		);
	END COMPONENT;
	--FOR ALL : busdr USE ENTITY work.busdr(one);

	COMPONENT reg16 IS
		PORT (
			din   : IN std_logic_vector(15 DOWNTO 0);
			dout  : OUT std_logic_vector(15 DOWNTO 0);
			load  : IN std_logic
		);
	END COMPONENT;
	--FOR ALL : reg16 USE ENTITY WORK.reg16(one);

	COMPONENT mux2_to_1x16 IS
		PORT (
			a, b    : IN std_logic_vector(15 DOWNTO 0);
			sa, sb  : IN std_logic;
			muxout  : OUT std_logic_vector(15 DOWNTO 0)
		);
	END COMPONENT;
	SIGNAL mux0_out, regOut : std_logic_vector(15 DOWNTO 0);
	SIGNAL regLoad, Abusdr_load, Bbusdr_load : std_logic;

	BEGIN
		mux0 : mux2_to_1x16
		PORT MAP(ABUS, BBUS, Arsel, Brsel, mux0_out);

		reg0 : reg16	PORT MAP(mux0_out, regOut, regLoad);
		Abusdr : busdr	PORT MAP(Abusdr_load, regOut, ABUS);
		Bbusdr : busdr	PORT MAP(Bbusdr_load, regOut, BBUS);

		Abusdr_load <= (Adrive) AND (Arsel);
		Bbusdr_load <= (Bdrive) AND (Brsel);
		regLoad <= (Aload AND Arsel) OR (Bload AND Brsel);
END one;