LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.std_logic_arith.ALL;
ENTITY tb4_1_MUX IS
END tb4_1_MUX;

ARCHITECTURE one OF tb4_1_MUX IS
	COMPONENT MUX_41_1_wide
		PORT (
			a, b, c, d, sel_0, sel_1  : IN std_logic;
			z                         : OUT std_logic
		);
	END COMPONENT;

	SIGNAL a, b, c, d, sel_0, sel_1, z : std_logic := '0';
	SIGNAL s1 : std_logic_vector(3 DOWNTO 0);
	SIGNAL i,j : INTEGER := 0;

	SIGNAL clk : BIT := '1';
BEGIN
	mux1 : MUX_41_1_wide PORT MAP(a, b, c, d, sel_0, sel_1, z);
 
 
	clk <= NOT clk AFTER 10 ns;
 
	PROCESS (clk)
	BEGIN
		IF (i < 16) THEN
			s1 <= conv_std_logic_vector(i, s1'length);
			a <= s1(0);
			b <= s1(1);
			c <= s1(2);
			d <= s1(3);
			i <= i + 1;
		ELSE
			i <= 0;
			j <= j + 1;
			sel_0 <= NOT sel_0;
		END IF;
		IF(j > 1 AND j < 4) THEN
		sel_1 <= '1';
		ELSE
		sel_1 <='0';
		END IF;

	END PROCESS;

END one;